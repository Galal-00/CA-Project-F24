LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

entity IF is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        -- Inputs
        
        
    );
end entity;